module bsg_iterative_cpa #(
  parameter integer width_p = 64
)